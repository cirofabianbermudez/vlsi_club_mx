module ROM_signal (
	
    input  LDX,  				// Toma siguiente valor
    output reg [15:0] DATTA  	// Datos de salida de 16 bits
);

    // Definir la ROM como una matriz de 200 palabras de 16 bits
    
	reg [7:0] addr=0;
	reg [15:0] rom [0:199];
	
	always @(*)	 begin
		if(LDX & addr < 200)
			addr = addr + 1;
			
		if ( addr == 200)
			addr = 0; 
		else
			addr <= addr;
			end

    initial begin
        rom[0] = 16'b0000000000000000;
        rom[1] = 16'b0000000011101110;
        rom[2] = 16'b1111111101100101;
        rom[3] = 16'b0000001010111100;
        rom[4] = 16'b1111111011011101;
        rom[5] = 16'b0000010001100100;
        rom[6] = 16'b1111111001111101;
        rom[7] = 16'b0000010111001110;
        rom[8] = 16'b1111111001010011;
        rom[9] = 16'b0000011011100111;
        rom[10] = 16'b1111111001101011;
        rom[11] = 16'b0000011110100011;
        rom[12] = 16'b1111111011001010;
        rom[13] = 16'b0000011111111010;
        rom[14] = 16'b1111111101101110;
        rom[15] = 16'b0000011111101011;
        rom[16] = 16'b0000000001010011;
        rom[17] = 16'b0000011101111110;
        rom[18] = 16'b0000000101101010;
        rom[19] = 16'b0000011010111101;
        rom[20] = 16'b0000001010100100;
        rom[21] = 16'b0000010110111011;
        rom[22] = 16'b0000001111101010;
        rom[23] = 16'b0000010010001100;
        rom[24] = 16'b0000010100100111;
        rom[25] = 16'b0000001101000111;
        rom[26] = 16'b0000011001000011;
        rom[27] = 16'b0000001000000100;
        rom[28] = 16'b0000011100100111;
        rom[29] = 16'b0000000011011001;
        rom[30] = 16'b0000011111000000;
        rom[31] = 16'b1111111111011001;
        rom[32] = 16'b0000011111111111;
        rom[33] = 16'b1111111100010011;
        rom[34] = 16'b0000011111011011;
        rom[35] = 16'b1111111010010001;
        rom[36] = 16'b0000011101010010;
        rom[37] = 16'b1111111001010111;
        rom[38] = 16'b0000011001100110;
        rom[39] = 16'b1111111001100001;
        rom[40] = 16'b0000010100100010;
        rom[41] = 16'b1111111010100111;
        rom[42] = 16'b0000001110010111;
        rom[43] = 16'b1111111100011101;
        rom[44] = 16'b0000000111011000;
        rom[45] = 16'b1111111110110001;
        rom[46] = 16'b0000000000000000;
        rom[47] = 16'b0000000001001111;
        rom[48] = 16'b1111111000101000;
        rom[49] = 16'b0000000011100011;
        rom[50] = 16'b1111110001101001;
        rom[51] = 16'b0000000101011001;
        rom[52] = 16'b1111101011011110;
        rom[53] = 16'b0000000110011111;
        rom[54] = 16'b1111100110011010;
        rom[55] = 16'b0000000110101001;
        rom[56] = 16'b1111100010101110;
        rom[57] = 16'b0000000101101111;
        rom[58] = 16'b1111100000100101;
        rom[59] = 16'b0000000011101101;
        rom[60] = 16'b1111100000000001;
        rom[61] = 16'b0000000000100111;
        rom[62] = 16'b1111100001000000;
        rom[63] = 16'b1111111100100111;
        rom[64] = 16'b1111100011011001;
        rom[65] = 16'b1111110111111100;
        rom[66] = 16'b1111100110111101;
        rom[67] = 16'b1111110010111001;
        rom[68] = 16'b1111101011011001;
        rom[69] = 16'b1111101101110100;
        rom[70] = 16'b1111110000010110;
        rom[71] = 16'b1111101001000101;
        rom[72] = 16'b1111110101011100;
        rom[73] = 16'b1111100101000011;
        rom[74] = 16'b1111111010010110;
        rom[75] = 16'b1111100010000010;
        rom[76] = 16'b1111111110101101;
        rom[77] = 16'b1111100000010101;
        rom[78] = 16'b0000000010010010;
        rom[79] = 16'b1111100000000110;
        rom[80] = 16'b0000000100110110;
        rom[81] = 16'b1111100001011101;
        rom[82] = 16'b0000000110010101;
        rom[83] = 16'b1111100100011001;
        rom[84] = 16'b0000000110101101;
        rom[85] = 16'b1111101000110010;
        rom[86] = 16'b0000000110000011;
        rom[87] = 16'b1111101110011100;
        rom[88] = 16'b0000000100100011;
        rom[89] = 16'b1111110101000100;
        rom[90] = 16'b0000000010011011;
        rom[91] = 16'b1111111100010010;
        rom[92] = 16'b0000000000000000;
        rom[93] = 16'b0000000011101110;
        rom[94] = 16'b1111111101100101;
        rom[95] = 16'b0000001010111100;
        rom[96] = 16'b1111111011011101;
        rom[97] = 16'b0000010001100100;
        rom[98] = 16'b1111111001111101;
        rom[99] = 16'b0000010111001110;
        rom[100] = 16'b1111111001010011;
        rom[101] = 16'b0000011011100111;
        rom[102] = 16'b1111111001101011;
        rom[103] = 16'b0000011110100011;
        rom[104] = 16'b1111111011001010;
        rom[105] = 16'b0000011111111010;
        rom[106] = 16'b1111111101101110;
        rom[107] = 16'b0000011111101011;
        rom[108] = 16'b0000000001010011;
        rom[109] = 16'b0000011101111110;
        rom[110] = 16'b0000000101101010;
        rom[111] = 16'b0000011010111101;
        rom[112] = 16'b0000001010100100;
        rom[113] = 16'b0000010110111011;
        rom[114] = 16'b0000001111101010;
        rom[115] = 16'b0000010010001100;
        rom[116] = 16'b0000010100100111;
        rom[117] = 16'b0000001101000111;
        rom[118] = 16'b0000011001000011;
        rom[119] = 16'b0000001000000100;
        rom[120] = 16'b0000011100100111;
        rom[121] = 16'b0000000011011001;
        rom[122] = 16'b0000011111000000;
        rom[123] = 16'b1111111111011001;
        rom[124] = 16'b0000011111111111;
        rom[125] = 16'b1111111100010011;
        rom[126] = 16'b0000011111011011;
        rom[127] = 16'b1111111010010001;
        rom[128] = 16'b0000011101010010;
        rom[129] = 16'b1111111001010111;
        rom[130] = 16'b0000011001100110;
        rom[131] = 16'b1111111001100001;
        rom[132] = 16'b0000010100100010;
        rom[133] = 16'b1111111010100111;
        rom[134] = 16'b0000001110010111;
        rom[135] = 16'b1111111100011101;
        rom[136] = 16'b0000000111011000;
        rom[137] = 16'b1111111110110001;
        rom[138] = 16'b0000000000000000;
        rom[139] = 16'b0000000001001111;
        rom[140] = 16'b1111111000101000;
        rom[141] = 16'b0000000011100011;
        rom[142] = 16'b1111110001101001;
        rom[143] = 16'b0000000101011001;
        rom[144] = 16'b1111101011011110;
        rom[145] = 16'b0000000110011111;
        rom[146] = 16'b1111100110011010;
        rom[147] = 16'b0000000110101001;
        rom[148] = 16'b1111100010101110;
        rom[149] = 16'b0000000101101111;
        rom[150] = 16'b1111100000100101;
        rom[151] = 16'b0000000011101101;
        rom[152] = 16'b1111100000000001;
        rom[153] = 16'b0000000000100111;
        rom[154] = 16'b1111100001000000;
        rom[155] = 16'b1111111100100111;
        rom[156] = 16'b1111100011011001;
        rom[157] = 16'b1111110111111100;
        rom[158] = 16'b1111100110111101;
        rom[159] = 16'b1111110010111001;
        rom[160] = 16'b1111101011011001;
        rom[161] = 16'b1111101101110100;
        rom[162] = 16'b1111110000010110;
        rom[163] = 16'b1111101001000101;
        rom[164] = 16'b1111110101011100;
        rom[165] = 16'b1111100101000011;
        rom[166] = 16'b1111111010010110;
        rom[167] = 16'b1111100010000010;
        rom[168] = 16'b1111111110101101;
        rom[169] = 16'b1111100000010101;
        rom[170] = 16'b0000000010010010;
        rom[171] = 16'b1111100000000110;
        rom[172] = 16'b0000000100110110;
        rom[173] = 16'b1111100001011101;
        rom[174] = 16'b0000000110010101;
        rom[175] = 16'b1111100100011001;
        rom[176] = 16'b0000000110101101;
        rom[177] = 16'b1111101000110010;
        rom[178] = 16'b0000000110000011;
        rom[179] = 16'b1111101110011100;
        rom[180] = 16'b0000000100100011;
        rom[181] = 16'b1111110101000100;
        rom[182] = 16'b0000000010011011;
        rom[183] = 16'b1111111100010010;
        rom[184] = 16'b0000000000000000;
        rom[185] = 16'b0000000011101110;
        rom[186] = 16'b1111111101100101;
        rom[187] = 16'b0000001010111100;
        rom[188] = 16'b1111111011011101;
        rom[189] = 16'b0000010001100100;
        rom[190] = 16'b1111111001111101;
        rom[191] = 16'b0000010111001110;
        rom[192] = 16'b1111111001010011;
        rom[193] = 16'b0000011011100111;
        rom[194] = 16'b1111111001101011;
        rom[195] = 16'b0000011110100011;
        rom[196] = 16'b1111111011001010;
        rom[197] = 16'b0000011111111010;
        rom[198] = 16'b1111111101101110;
        rom[199] = 16'b0000011111101011;
    end

    // Asignar el valor de la ROM a la salida en base a la direcci n
    always @(*) begin
        DATTA = rom[addr];
    end

endmodule
